/*
 * Tiny Canvas - MS Paint Style Drawing Tool
 * Gamepad-controlled pixel art with brush sizes, symmetry, and shapes.
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,
    output wire [7:0] uo_out,
    input  wire [7:0] uio_in,
    output wire [7:0] uio_out,
    output wire [7:0] uio_oe,
    input  wire       ena,
    input  wire       clk,
    input  wire       rst_n
);

    // ================================================================
    // Gamepad PMOD Input
    // ================================================================
    wire pmod_data  = ui_in[0];
    wire pmod_clk   = ui_in[1];
    wire pmod_latch = ui_in[2];

    wire gp_b, gp_y, gp_select, gp_start;
    wire gp_up, gp_down, gp_left, gp_right;
    wire gp_a, gp_x, gp_l, gp_r;
    wire gp_is_present;

    gamepad_pmod_single gamepad_inst (
        .rst_n(rst_n), .clk(clk),
        .pmod_data(pmod_data), .pmod_clk(pmod_clk), .pmod_latch(pmod_latch),
        .b(gp_b), .y(gp_y), .select(gp_select), .start(gp_start),
        .up(gp_up), .down(gp_down), .left(gp_left), .right(gp_right),
        .a(gp_a), .x(gp_x), .l(gp_l), .r(gp_r),
        .is_present(gp_is_present)
    );

    // ================================================================
    // Button Edge Detection & Toggle Logic
    // ================================================================
    reg y_prev, x_prev, b_prev, a_prev;
    reg sw_red, sw_green, sw_blue, brush_mode;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            y_prev <= 1'b0; x_prev <= 1'b0; b_prev <= 1'b0; a_prev <= 1'b0;
            sw_red <= 1'b0; sw_green <= 1'b0; sw_blue <= 1'b0;
            brush_mode <= 1'b1;
        end else begin
            y_prev <= gp_y; x_prev <= gp_x; b_prev <= gp_b; a_prev <= gp_a;
            
            if (gp_y && !y_prev) sw_red <= ~sw_red;
            if (gp_x && !x_prev) sw_green <= ~sw_green;
            if (gp_b && !b_prev) sw_blue <= ~sw_blue;
            if (gp_a && !a_prev) brush_mode <= ~brush_mode;
        end
    end

    // ================================================================
    // Position Tracker
    // ================================================================
    wire [7:0] x_pos, y_pos;
    wire [3:0] dir_udlr = {gp_up, gp_down, gp_left, gp_right};
    wire movement = gp_up || gp_down || gp_left || gp_right;
    reg movement_prev;
    wire movement_edge = movement && !movement_prev;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) movement_prev <= 1'b0;
        else movement_prev <= movement;
    end

    position pos_inst (
        .x_pos(x_pos), .y_pos(y_pos),
        .dir_udlr(dir_udlr),
        .clk(clk), .rst_n(rst_n)
    );

    // ================================================================
    // Colour Mixing
    // ================================================================
    wire [2:0] colour_out;
    wire paint_enable;

    colour colour_inst (
        .clk(clk), .rst_n(rst_n),
        .sw_red(sw_red), .sw_green(sw_green), .sw_blue(sw_blue),
        .brush_mode(brush_mode),
        .colour_out(colour_out),
        .paint_enable(paint_enable)
    );

    // ================================================================
    // Brush Settings (L/R = size, Start = symmetry)
    // ================================================================
    wire [2:0] brush_size;
    wire [1:0] symmetry_mode;

    brush_settings brush_inst (
        .clk(clk), .rst_n(rst_n),
        .btn_size_up(gp_r),
        .btn_size_down(gp_l),
        .btn_symmetry(gp_start),
        .brush_size(brush_size),
        .symmetry_mode(symmetry_mode)
    );

    // ================================================================
    // Draw Mode (Select = cycle mode, A = set point)
    // ================================================================
    wire [1:0] draw_mode_out;
    wire [7:0] point_a_x, point_a_y, point_b_x, point_b_y;
    wire point_a_valid, shape_trigger;

    draw_mode mode_inst (
        .clk(clk), .rst_n(rst_n),
        .btn_mode(gp_select),
        .btn_point(gp_a),
        .x_pos(x_pos), .y_pos(y_pos),
        .mode(draw_mode_out),
        .point_a_x(point_a_x), .point_a_y(point_a_y),
        .point_a_valid(point_a_valid),
        .point_b_x(point_b_x), .point_b_y(point_b_y),
        .shape_trigger(shape_trigger)
    );

    // ================================================================
    // Draw Engine (coordinates freehand, line, rect, spray)
    // ================================================================
    wire [7:0] draw_x, draw_y;
    wire draw_valid, draw_busy;

    draw_engine engine_inst (
        .clk(clk), .rst_n(rst_n),
        .mode(draw_mode_out),
        .x_pos(x_pos), .y_pos(y_pos),
        .move_trigger(movement_edge),
        .shape_trigger(shape_trigger),
        .point_a_x(point_a_x), .point_a_y(point_a_y),
        .point_b_x(point_b_x), .point_b_y(point_b_y),
        .paint_enable(paint_enable),
        .pixel_x(draw_x), .pixel_y(draw_y),
        .pixel_valid(draw_valid),
        .busy(draw_busy)
    );

    // ================================================================
    // Packet Generator (expands brush size + symmetry)
    // ================================================================
    wire [7:0] pkt_x, pkt_y;
    wire pkt_valid, pkt_busy;

    packet_generator pkt_inst (
        .clk(clk), .rst_n(rst_n),
        .trigger(draw_valid),
        .x_in(draw_x), .y_in(draw_y),
        .brush_size(brush_size),
        .symmetry_mode(symmetry_mode),
        .x_out(pkt_x), .y_out(pkt_y),
        .valid(pkt_valid),
        .busy(pkt_busy)
    );

    // ================================================================
    // Status Byte Construction
    // ================================================================
    wire [7:0] status_reg;
    assign status_reg[7]   = gp_up;
    assign status_reg[6]   = gp_down;
    assign status_reg[5]   = gp_left;
    assign status_reg[4]   = gp_right;
    assign status_reg[3]   = brush_mode;
    assign status_reg[2:0] = colour_out;

    // ================================================================
    // I2C Slave Interface
    // ================================================================
    wire sda_oe_int, sda_out_int;

    i2c_slave #(.I2C_ADDR(7'b1100100)) i2c_slave_inst (
        .scl(uio_in[2]),
        .sda_in(uio_in[1]),
        .sda_oe(sda_oe_int),
        .sda_out(sda_out_int),
        .i2c_state(uo_out[2:0]),
        .x_pos(pkt_x),
        .y_pos(pkt_y),
        .status(status_reg),
        .clk(clk),
        .rst_n(rst_n)
    );

    // ================================================================
    // I/O Wiring
    // ================================================================
    assign uio_out[1] = 1'b0;
    assign uio_oe[1]  = sda_oe_int;
    assign uio_out[2] = 1'b0;
    assign uio_oe[2]  = 1'b0;
    assign uio_out[7:3] = 5'b0;
    assign uio_oe[7:3]  = 5'b0;
    assign uio_out[0]   = 1'b0;
    assign uio_oe[0]    = 1'b0;
    assign uo_out[7:3] = 5'b0;

    // ================================================================
    // Unused Signals
    // ================================================================
    wire _unused = &{ena, sda_out_int, ui_in[7:3], uio_in[7:3], uio_in[0],
                     gp_is_present, draw_busy, pkt_busy, point_a_valid};

endmodule
